module top (
    input  wire         clk,
    input  wire         rstn);

    cpu(clk, rstn);

endmodule

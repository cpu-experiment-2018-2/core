interface gpr_if;
    reg signed [31:0] gpr [0:31];
endinterface
